module ALUcontrol(
  input  [2:0] io_aluOP,
  input  [2:0] io_fun_3,
  input        io_fun_7,
  output [4:0] io_aluControl
);
  wire  _T; // @[ALUcontrol.scala 16:20]
  wire  _T_1; // @[ALUcontrol.scala 16:40]
  wire  _T_2; // @[ALUcontrol.scala 16:28]
  wire [3:0] _T_3; // @[Cat.scala 29:58]
  wire  _T_6; // @[ALUcontrol.scala 19:33]
  wire [3:0] _T_7; // @[Cat.scala 29:58]
  wire  _T_8; // @[ALUcontrol.scala 22:25]
  wire  _T_9; // @[ALUcontrol.scala 22:45]
  wire  _T_10; // @[ALUcontrol.scala 22:33]
  wire  _T_12; // @[ALUcontrol.scala 22:53]
  wire  _T_18; // @[ALUcontrol.scala 25:53]
  wire  _T_21; // @[ALUcontrol.scala 28:45]
  wire  _T_22; // @[ALUcontrol.scala 28:33]
  wire  _T_26; // @[ALUcontrol.scala 34:25]
  wire [4:0] _T_27; // @[Cat.scala 29:58]
  wire  _T_28; // @[ALUcontrol.scala 37:25]
  wire [4:0] _GEN_0; // @[ALUcontrol.scala 37:33]
  wire [4:0] _GEN_1; // @[ALUcontrol.scala 34:33]
  wire [4:0] _GEN_2; // @[ALUcontrol.scala 31:33]
  wire [4:0] _GEN_3; // @[ALUcontrol.scala 28:53]
  wire [4:0] _GEN_4; // @[ALUcontrol.scala 25:73]
  wire [4:0] _GEN_5; // @[ALUcontrol.scala 22:73]
  wire [4:0] _GEN_6; // @[ALUcontrol.scala 19:53]
  assign _T = io_aluOP == 3'h0; // @[ALUcontrol.scala 16:20]
  assign _T_1 = io_fun_7 == 1'h0; // @[ALUcontrol.scala 16:40]
  assign _T_2 = _T & _T_1; // @[ALUcontrol.scala 16:28]
  assign _T_3 = {1'h0,io_fun_3}; // @[Cat.scala 29:58]
  assign _T_6 = _T & io_fun_7; // @[ALUcontrol.scala 19:33]
  assign _T_7 = {1'h1,io_fun_3}; // @[Cat.scala 29:58]
  assign _T_8 = io_aluOP == 3'h1; // @[ALUcontrol.scala 22:25]
  assign _T_9 = io_fun_3 == 3'h5; // @[ALUcontrol.scala 22:45]
  assign _T_10 = _T_8 & _T_9; // @[ALUcontrol.scala 22:33]
  assign _T_12 = _T_10 & _T_1; // @[ALUcontrol.scala 22:53]
  assign _T_18 = _T_10 & io_fun_7; // @[ALUcontrol.scala 25:53]
  assign _T_21 = io_fun_3 == 3'h1; // @[ALUcontrol.scala 28:45]
  assign _T_22 = _T_8 & _T_21; // @[ALUcontrol.scala 28:33]
  assign _T_26 = io_aluOP == 3'h2; // @[ALUcontrol.scala 34:25]
  assign _T_27 = {2'h2,io_fun_3}; // @[Cat.scala 29:58]
  assign _T_28 = io_aluOP == 3'h3; // @[ALUcontrol.scala 37:25]
  assign _GEN_0 = _T_28 ? 5'h1f : 5'h0; // @[ALUcontrol.scala 37:33]
  assign _GEN_1 = _T_26 ? _T_27 : _GEN_0; // @[ALUcontrol.scala 34:33]
  assign _GEN_2 = _T_8 ? {{1'd0}, _T_3} : _GEN_1; // @[ALUcontrol.scala 31:33]
  assign _GEN_3 = _T_22 ? {{1'd0}, _T_3} : _GEN_2; // @[ALUcontrol.scala 28:53]
  assign _GEN_4 = _T_18 ? {{1'd0}, _T_7} : _GEN_3; // @[ALUcontrol.scala 25:73]
  assign _GEN_5 = _T_12 ? {{1'd0}, _T_3} : _GEN_4; // @[ALUcontrol.scala 22:73]
  assign _GEN_6 = _T_6 ? {{1'd0}, _T_7} : _GEN_5; // @[ALUcontrol.scala 19:53]
  assign io_aluControl = _T_2 ? {{1'd0}, _T_3} : _GEN_6; // @[ALUcontrol.scala 14:19 ALUcontrol.scala 17:23 ALUcontrol.scala 20:23 ALUcontrol.scala 23:23 ALUcontrol.scala 26:23 ALUcontrol.scala 29:23 ALUcontrol.scala 32:23 ALUcontrol.scala 35:23 ALUcontrol.scala 38:23 ALUcontrol.scala 41:23]
endmodule