module ALU(
  input  [31:0] io_oprndA,
  input  [31:0] io_oprndB,
  input  [4:0]  io_aluControl,
  output        io_branch,
  output [31:0] io_aluOUT
);
  wire [4:0] shamt; // @[ALU.scala 16:26]
  wire [1:0] _T; // @[ALU.scala 18:33]
  wire  _T_1; // @[ALU.scala 18:39]
  wire  _T_2; // @[ALU.scala 18:61]
  wire  _T_4; // @[ALU.scala 21:25]
  wire [31:0] _T_6; // @[ALU.scala 22:32]
  wire [31:0] _T_7; // @[ALU.scala 22:32]
  wire  _T_8; // @[ALU.scala 24:30]
  wire [62:0] _GEN_25; // @[ALU.scala 25:32]
  wire [62:0] _T_9; // @[ALU.scala 25:32]
  wire  _T_10; // @[ALU.scala 27:30]
  wire  _T_11; // @[ALU.scala 28:24]
  wire  _T_12; // @[ALU.scala 34:30]
  wire [31:0] _T_13; // @[ALU.scala 35:26]
  wire [31:0] _T_14; // @[ALU.scala 35:47]
  wire  _T_15; // @[ALU.scala 35:33]
  wire  _T_16; // @[ALU.scala 41:30]
  wire [31:0] _T_17; // @[ALU.scala 42:32]
  wire [31:0] _T_18; // @[ALU.scala 42:32]
  wire  _T_19; // @[ALU.scala 44:30]
  wire [31:0] _T_20; // @[ALU.scala 45:32]
  wire  _T_21; // @[ALU.scala 47:30]
  wire [31:0] _T_22; // @[ALU.scala 48:32]
  wire [31:0] _T_23; // @[ALU.scala 48:32]
  wire  _T_24; // @[ALU.scala 50:30]
  wire [31:0] _T_25; // @[ALU.scala 51:32]
  wire [31:0] _T_26; // @[ALU.scala 51:32]
  wire  _T_27; // @[ALU.scala 53:30]
  wire [31:0] _T_29; // @[ALU.scala 54:32]
  wire [31:0] _T_30; // @[ALU.scala 54:32]
  wire  _T_31; // @[ALU.scala 56:30]
  wire  _T_33; // @[ALU.scala 59:30]
  wire  _T_34; // @[ALU.scala 60:24]
  wire [1:0] _GEN_2; // @[ALU.scala 60:38]
  wire  _T_35; // @[ALU.scala 66:30]
  wire  _T_36; // @[ALU.scala 67:26]
  wire [1:0] _GEN_3; // @[ALU.scala 67:40]
  wire  _T_37; // @[ALU.scala 74:30]
  wire [1:0] _GEN_4; // @[ALU.scala 75:36]
  wire  _T_39; // @[ALU.scala 82:30]
  wire  _T_40; // @[ALU.scala 83:24]
  wire [1:0] _GEN_5; // @[ALU.scala 83:37]
  wire  _T_41; // @[ALU.scala 90:30]
  wire [1:0] _GEN_6; // @[ALU.scala 91:54]
  wire  _T_45; // @[ALU.scala 97:30]
  wire  _T_48; // @[ALU.scala 98:33]
  wire [1:0] _GEN_7; // @[ALU.scala 98:55]
  wire  _T_49; // @[ALU.scala 104:30]
  wire [31:0] _GEN_8; // @[ALU.scala 104:39]
  wire [31:0] _GEN_9; // @[ALU.scala 97:39]
  wire [31:0] _GEN_10; // @[ALU.scala 90:39]
  wire [31:0] _GEN_11; // @[ALU.scala 82:39]
  wire [31:0] _GEN_12; // @[ALU.scala 74:39]
  wire [31:0] _GEN_13; // @[ALU.scala 66:39]
  wire [31:0] _GEN_14; // @[ALU.scala 59:39]
  wire [31:0] _GEN_15; // @[ALU.scala 56:39]
  wire [31:0] _GEN_16; // @[ALU.scala 53:38]
  wire [31:0] _GEN_17; // @[ALU.scala 50:38]
  wire [31:0] _GEN_18; // @[ALU.scala 47:38]
  wire [31:0] _GEN_19; // @[ALU.scala 44:38]
  wire [31:0] _GEN_20; // @[ALU.scala 41:38]
  wire [31:0] _GEN_21; // @[ALU.scala 34:38]
  wire [31:0] _GEN_22; // @[ALU.scala 27:38]
  wire [62:0] _GEN_23; // @[ALU.scala 24:38]
  wire [62:0] _GEN_24; // @[ALU.scala 21:33]
  wire [31:0] _GEN_26; // @[ALU.scala 14:15 ALU.scala 22:19 ALU.scala 25:19 ALU.scala 29:23 ALU.scala 31:23 ALU.scala 36:23 ALU.scala 38:23 ALU.scala 42:19 ALU.scala 45:19 ALU.scala 48:19 ALU.scala 51:19 ALU.scala 54:19 ALU.scala 57:19 ALU.scala 61:23 ALU.scala 63:23 ALU.scala 68:25 ALU.scala 70:25 ALU.scala 76:23 ALU.scala 78:23 ALU.scala 84:23 ALU.scala 86:23 ALU.scala 92:23 ALU.scala 94:23 ALU.scala 99:23 ALU.scala 101:23 ALU.scala 105:19]
  assign shamt = io_oprndB[4:0]; // @[ALU.scala 16:26]
  assign _T = io_aluControl[4:3]; // @[ALU.scala 18:33]
  assign _T_1 = _T == 2'h2; // @[ALU.scala 18:39]
  assign _T_2 = $signed(io_aluOUT) == $signed(32'sh1); // @[ALU.scala 18:61]
  assign _T_4 = io_aluControl == 5'h0; // @[ALU.scala 21:25]
  assign _T_6 = $signed(io_oprndA) + $signed(io_oprndB); // @[ALU.scala 22:32]
  assign _T_7 = $signed(_T_6); // @[ALU.scala 22:32]
  assign _T_8 = io_aluControl == 5'h1; // @[ALU.scala 24:30]
  assign _GEN_25 = {{31{io_oprndA[31]}},io_oprndA}; // @[ALU.scala 25:32]
  assign _T_9 = $signed(_GEN_25) << shamt; // @[ALU.scala 25:32]
  assign _T_10 = io_aluControl == 5'h2; // @[ALU.scala 27:30]
  assign _T_11 = $signed(io_oprndA) < $signed(io_oprndB); // @[ALU.scala 28:24]
  assign _T_12 = io_aluControl == 5'h3; // @[ALU.scala 34:30]
  assign _T_13 = $unsigned(io_oprndA); // @[ALU.scala 35:26]
  assign _T_14 = $unsigned(io_oprndB); // @[ALU.scala 35:47]
  assign _T_15 = _T_13 < _T_14; // @[ALU.scala 35:33]
  assign _T_16 = io_aluControl == 5'h4; // @[ALU.scala 41:30]
  assign _T_17 = $signed(io_oprndA) ^ $signed(io_oprndB); // @[ALU.scala 42:32]
  assign _T_18 = $signed(_T_17); // @[ALU.scala 42:32]
  assign _T_19 = io_aluControl == 5'h5; // @[ALU.scala 44:30]
  assign _T_20 = $signed(io_oprndA) >>> shamt; // @[ALU.scala 45:32]
  assign _T_21 = io_aluControl == 5'h6; // @[ALU.scala 47:30]
  assign _T_22 = $signed(io_oprndA) | $signed(io_oprndB); // @[ALU.scala 48:32]
  assign _T_23 = $signed(_T_22); // @[ALU.scala 48:32]
  assign _T_24 = io_aluControl == 5'h7; // @[ALU.scala 50:30]
  assign _T_25 = $signed(io_oprndA) & $signed(io_oprndB); // @[ALU.scala 51:32]
  assign _T_26 = $signed(_T_25); // @[ALU.scala 51:32]
  assign _T_27 = io_aluControl == 5'h8; // @[ALU.scala 53:30]
  assign _T_29 = $signed(io_oprndA) - $signed(io_oprndB); // @[ALU.scala 54:32]
  assign _T_30 = $signed(_T_29); // @[ALU.scala 54:32]
  assign _T_31 = io_aluControl == 5'hd; // @[ALU.scala 56:30]
  assign _T_33 = io_aluControl == 5'h10; // @[ALU.scala 59:30]
  assign _T_34 = $signed(io_oprndA) == $signed(io_oprndB); // @[ALU.scala 60:24]
  assign _GEN_2 = _T_34 ? $signed(2'sh1) : $signed(2'sh0); // @[ALU.scala 60:38]
  assign _T_35 = io_aluControl == 5'h11; // @[ALU.scala 66:30]
  assign _T_36 = $signed(io_oprndA) != $signed(io_oprndB); // @[ALU.scala 67:26]
  assign _GEN_3 = _T_36 ? $signed(2'sh1) : $signed(2'sh0); // @[ALU.scala 67:40]
  assign _T_37 = io_aluControl == 5'h12; // @[ALU.scala 74:30]
  assign _GEN_4 = _T_11 ? $signed(2'sh1) : $signed(2'sh0); // @[ALU.scala 75:36]
  assign _T_39 = io_aluControl == 5'h13; // @[ALU.scala 82:30]
  assign _T_40 = $signed(io_oprndA) >= $signed(io_oprndB); // @[ALU.scala 83:24]
  assign _GEN_5 = _T_40 ? $signed(2'sh1) : $signed(2'sh0); // @[ALU.scala 83:37]
  assign _T_41 = io_aluControl == 5'h14; // @[ALU.scala 90:30]
  assign _GEN_6 = _T_15 ? $signed(2'sh1) : $signed(2'sh0); // @[ALU.scala 91:54]
  assign _T_45 = io_aluControl == 5'h15; // @[ALU.scala 97:30]
  assign _T_48 = _T_13 >= _T_14; // @[ALU.scala 98:33]
  assign _GEN_7 = _T_48 ? $signed(2'sh1) : $signed(2'sh0); // @[ALU.scala 98:55]
  assign _T_49 = io_aluControl == 5'h1f; // @[ALU.scala 104:30]
  assign _GEN_8 = _T_49 ? $signed(io_oprndA) : $signed(32'sh0); // @[ALU.scala 104:39]
  assign _GEN_9 = _T_45 ? $signed({{30{_GEN_7[1]}},_GEN_7}) : $signed(_GEN_8); // @[ALU.scala 97:39]
  assign _GEN_10 = _T_41 ? $signed({{30{_GEN_6[1]}},_GEN_6}) : $signed(_GEN_9); // @[ALU.scala 90:39]
  assign _GEN_11 = _T_39 ? $signed({{30{_GEN_5[1]}},_GEN_5}) : $signed(_GEN_10); // @[ALU.scala 82:39]
  assign _GEN_12 = _T_37 ? $signed({{30{_GEN_4[1]}},_GEN_4}) : $signed(_GEN_11); // @[ALU.scala 74:39]
  assign _GEN_13 = _T_35 ? $signed({{30{_GEN_3[1]}},_GEN_3}) : $signed(_GEN_12); // @[ALU.scala 66:39]
  assign _GEN_14 = _T_33 ? $signed({{30{_GEN_2[1]}},_GEN_2}) : $signed(_GEN_13); // @[ALU.scala 59:39]
  assign _GEN_15 = _T_31 ? $signed(_T_20) : $signed(_GEN_14); // @[ALU.scala 56:39]
  assign _GEN_16 = _T_27 ? $signed(_T_30) : $signed(_GEN_15); // @[ALU.scala 53:38]
  assign _GEN_17 = _T_24 ? $signed(_T_26) : $signed(_GEN_16); // @[ALU.scala 50:38]
  assign _GEN_18 = _T_21 ? $signed(_T_23) : $signed(_GEN_17); // @[ALU.scala 47:38]
  assign _GEN_19 = _T_19 ? $signed(_T_20) : $signed(_GEN_18); // @[ALU.scala 44:38]
  assign _GEN_20 = _T_16 ? $signed(_T_18) : $signed(_GEN_19); // @[ALU.scala 41:38]
  assign _GEN_21 = _T_12 ? $signed(32'sh1) : $signed(_GEN_20); // @[ALU.scala 34:38]
  assign _GEN_22 = _T_10 ? $signed(32'sh1) : $signed(_GEN_21); // @[ALU.scala 27:38]
  assign _GEN_23 = _T_8 ? $signed(_T_9) : $signed({{31{_GEN_22[31]}},_GEN_22}); // @[ALU.scala 24:38]
  assign _GEN_24 = _T_4 ? $signed({{31{_T_7[31]}},_T_7}) : $signed(_GEN_23); // @[ALU.scala 21:33]
  assign io_branch = _T_1 & _T_2; // @[ALU.scala 18:15]
  assign _GEN_26 = _GEN_24[31:0]; // @[ALU.scala 14:15 ALU.scala 22:19 ALU.scala 25:19 ALU.scala 29:23 ALU.scala 31:23 ALU.scala 36:23 ALU.scala 38:23 ALU.scala 42:19 ALU.scala 45:19 ALU.scala 48:19 ALU.scala 51:19 ALU.scala 54:19 ALU.scala 57:19 ALU.scala 61:23 ALU.scala 63:23 ALU.scala 68:25 ALU.scala 70:25 ALU.scala 76:23 ALU.scala 78:23 ALU.scala 84:23 ALU.scala 86:23 ALU.scala 92:23 ALU.scala 94:23 ALU.scala 99:23 ALU.scala 101:23 ALU.scala 105:19]
  assign io_aluOUT = $signed(_GEN_26); // @[ALU.scala 14:15 ALU.scala 22:19 ALU.scala 25:19 ALU.scala 29:23 ALU.scala 31:23 ALU.scala 36:23 ALU.scala 38:23 ALU.scala 42:19 ALU.scala 45:19 ALU.scala 48:19 ALU.scala 51:19 ALU.scala 54:19 ALU.scala 57:19 ALU.scala 61:23 ALU.scala 63:23 ALU.scala 68:25 ALU.scala 70:25 ALU.scala 76:23 ALU.scala 78:23 ALU.scala 84:23 ALU.scala 86:23 ALU.scala 92:23 ALU.scala 94:23 ALU.scala 99:23 ALU.scala 101:23 ALU.scala 105:19]
endmodule