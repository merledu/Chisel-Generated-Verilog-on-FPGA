module ControlDecode(
  input        io_rtype,
  input        io_itype,
  input        io_load,
  input        io_stype,
  input        io_sbtype,
  input        io_lui,
  input        io_auipc,
  input        io_ujtype,
  input        io_jalr,
  output       io_regWrite,
  output       io_memtoReg,
  output       io_memRead,
  output       io_memWrite,
  output       io_branch,
  output [1:0] io_oprndAsel,
  output       io_oprndBsel,
  output [1:0] io_immSel,
  output [1:0] io_nextPCsel,
  output [2:0] io_aluOP
);
  wire [1:0] _GEN_1; // @[ControlDecode.scala 84:28]
  wire [1:0] _GEN_2; // @[ControlDecode.scala 84:28]
  wire  _GEN_3; // @[ControlDecode.scala 78:30]
  wire [1:0] _GEN_4; // @[ControlDecode.scala 78:30]
  wire [1:0] _GEN_5; // @[ControlDecode.scala 78:30]
  wire [1:0] _GEN_6; // @[ControlDecode.scala 78:30]
  wire  _GEN_7; // @[ControlDecode.scala 71:29]
  wire [1:0] _GEN_8; // @[ControlDecode.scala 71:29]
  wire [1:0] _GEN_10; // @[ControlDecode.scala 71:29]
  wire [2:0] _GEN_11; // @[ControlDecode.scala 71:29]
  wire [1:0] _GEN_12; // @[ControlDecode.scala 71:29]
  wire  _GEN_13; // @[ControlDecode.scala 65:27]
  wire  _GEN_14; // @[ControlDecode.scala 65:27]
  wire [1:0] _GEN_15; // @[ControlDecode.scala 65:27]
  wire [2:0] _GEN_16; // @[ControlDecode.scala 65:27]
  wire [1:0] _GEN_17; // @[ControlDecode.scala 65:27]
  wire [1:0] _GEN_18; // @[ControlDecode.scala 65:27]
  wire [1:0] _GEN_20; // @[ControlDecode.scala 60:30]
  wire [2:0] _GEN_21; // @[ControlDecode.scala 60:30]
  wire  _GEN_22; // @[ControlDecode.scala 60:30]
  wire  _GEN_23; // @[ControlDecode.scala 60:30]
  wire [1:0] _GEN_24; // @[ControlDecode.scala 60:30]
  wire [1:0] _GEN_25; // @[ControlDecode.scala 60:30]
  wire  _GEN_27; // @[ControlDecode.scala 54:29]
  wire [1:0] _GEN_28; // @[ControlDecode.scala 54:29]
  wire [2:0] _GEN_29; // @[ControlDecode.scala 54:29]
  wire  _GEN_30; // @[ControlDecode.scala 54:29]
  wire [1:0] _GEN_31; // @[ControlDecode.scala 54:29]
  wire  _GEN_32; // @[ControlDecode.scala 54:29]
  wire [1:0] _GEN_33; // @[ControlDecode.scala 54:29]
  wire  _GEN_34; // @[ControlDecode.scala 47:28]
  wire  _GEN_36; // @[ControlDecode.scala 47:28]
  wire [2:0] _GEN_37; // @[ControlDecode.scala 47:28]
  wire  _GEN_38; // @[ControlDecode.scala 47:28]
  wire [1:0] _GEN_39; // @[ControlDecode.scala 47:28]
  wire  _GEN_40; // @[ControlDecode.scala 47:28]
  wire [1:0] _GEN_41; // @[ControlDecode.scala 47:28]
  wire [1:0] _GEN_42; // @[ControlDecode.scala 47:28]
  wire  _GEN_43; // @[ControlDecode.scala 42:29]
  wire  _GEN_44; // @[ControlDecode.scala 42:29]
  wire [2:0] _GEN_45; // @[ControlDecode.scala 42:29]
  wire  _GEN_46; // @[ControlDecode.scala 42:29]
  wire  _GEN_47; // @[ControlDecode.scala 42:29]
  wire [1:0] _GEN_48; // @[ControlDecode.scala 42:29]
  wire  _GEN_49; // @[ControlDecode.scala 42:29]
  wire [1:0] _GEN_50; // @[ControlDecode.scala 42:29]
  wire [1:0] _GEN_51; // @[ControlDecode.scala 42:29]
  assign _GEN_1 = io_jalr ? 2'h2 : 2'h0; // @[ControlDecode.scala 84:28]
  assign _GEN_2 = io_jalr ? 2'h3 : 2'h0; // @[ControlDecode.scala 84:28]
  assign _GEN_3 = io_ujtype | io_jalr; // @[ControlDecode.scala 78:30]
  assign _GEN_4 = io_ujtype ? 2'h2 : _GEN_1; // @[ControlDecode.scala 78:30]
  assign _GEN_5 = io_ujtype ? 2'h2 : _GEN_2; // @[ControlDecode.scala 78:30]
  assign _GEN_6 = io_ujtype ? 2'h3 : _GEN_2; // @[ControlDecode.scala 78:30]
  assign _GEN_7 = io_auipc | _GEN_3; // @[ControlDecode.scala 71:29]
  assign _GEN_8 = io_auipc ? 2'h1 : _GEN_4; // @[ControlDecode.scala 71:29]
  assign _GEN_10 = io_auipc ? 2'h2 : 2'h0; // @[ControlDecode.scala 71:29]
  assign _GEN_11 = io_auipc ? 3'h4 : {{1'd0}, _GEN_6}; // @[ControlDecode.scala 71:29]
  assign _GEN_12 = io_auipc ? 2'h0 : _GEN_5; // @[ControlDecode.scala 71:29]
  assign _GEN_13 = io_lui | _GEN_7; // @[ControlDecode.scala 65:27]
  assign _GEN_14 = io_lui | io_auipc; // @[ControlDecode.scala 65:27]
  assign _GEN_15 = io_lui ? 2'h2 : _GEN_10; // @[ControlDecode.scala 65:27]
  assign _GEN_16 = io_lui ? 3'h4 : _GEN_11; // @[ControlDecode.scala 65:27]
  assign _GEN_17 = io_lui ? 2'h0 : _GEN_8; // @[ControlDecode.scala 65:27]
  assign _GEN_18 = io_lui ? 2'h0 : _GEN_12; // @[ControlDecode.scala 65:27]
  assign _GEN_20 = io_sbtype ? 2'h1 : _GEN_18; // @[ControlDecode.scala 60:30]
  assign _GEN_21 = io_sbtype ? 3'h2 : _GEN_16; // @[ControlDecode.scala 60:30]
  assign _GEN_22 = io_sbtype ? 1'h0 : _GEN_13; // @[ControlDecode.scala 60:30]
  assign _GEN_23 = io_sbtype ? 1'h0 : _GEN_14; // @[ControlDecode.scala 60:30]
  assign _GEN_24 = io_sbtype ? 2'h0 : _GEN_15; // @[ControlDecode.scala 60:30]
  assign _GEN_25 = io_sbtype ? 2'h0 : _GEN_17; // @[ControlDecode.scala 60:30]
  assign _GEN_27 = io_stype | _GEN_23; // @[ControlDecode.scala 54:29]
  assign _GEN_28 = io_stype ? 2'h1 : _GEN_24; // @[ControlDecode.scala 54:29]
  assign _GEN_29 = io_stype ? 3'h4 : _GEN_21; // @[ControlDecode.scala 54:29]
  assign _GEN_30 = io_stype ? 1'h0 : io_sbtype; // @[ControlDecode.scala 54:29]
  assign _GEN_31 = io_stype ? 2'h0 : _GEN_20; // @[ControlDecode.scala 54:29]
  assign _GEN_32 = io_stype ? 1'h0 : _GEN_22; // @[ControlDecode.scala 54:29]
  assign _GEN_33 = io_stype ? 2'h0 : _GEN_25; // @[ControlDecode.scala 54:29]
  assign _GEN_34 = io_load | _GEN_32; // @[ControlDecode.scala 47:28]
  assign _GEN_36 = io_load | _GEN_27; // @[ControlDecode.scala 47:28]
  assign _GEN_37 = io_load ? 3'h4 : _GEN_29; // @[ControlDecode.scala 47:28]
  assign _GEN_38 = io_load ? 1'h0 : io_stype; // @[ControlDecode.scala 47:28]
  assign _GEN_39 = io_load ? 2'h0 : _GEN_28; // @[ControlDecode.scala 47:28]
  assign _GEN_40 = io_load ? 1'h0 : _GEN_30; // @[ControlDecode.scala 47:28]
  assign _GEN_41 = io_load ? 2'h0 : _GEN_31; // @[ControlDecode.scala 47:28]
  assign _GEN_42 = io_load ? 2'h0 : _GEN_33; // @[ControlDecode.scala 47:28]
  assign _GEN_43 = io_itype | _GEN_34; // @[ControlDecode.scala 42:29]
  assign _GEN_44 = io_itype | _GEN_36; // @[ControlDecode.scala 42:29]
  assign _GEN_45 = io_itype ? 3'h1 : _GEN_37; // @[ControlDecode.scala 42:29]
  assign _GEN_46 = io_itype ? 1'h0 : io_load; // @[ControlDecode.scala 42:29]
  assign _GEN_47 = io_itype ? 1'h0 : _GEN_38; // @[ControlDecode.scala 42:29]
  assign _GEN_48 = io_itype ? 2'h0 : _GEN_39; // @[ControlDecode.scala 42:29]
  assign _GEN_49 = io_itype ? 1'h0 : _GEN_40; // @[ControlDecode.scala 42:29]
  assign _GEN_50 = io_itype ? 2'h0 : _GEN_41; // @[ControlDecode.scala 42:29]
  assign _GEN_51 = io_itype ? 2'h0 : _GEN_42; // @[ControlDecode.scala 42:29]
  assign io_regWrite = io_rtype | _GEN_43; // @[ControlDecode.scala 28:17 ControlDecode.scala 40:17 ControlDecode.scala 43:17 ControlDecode.scala 48:17 ControlDecode.scala 66:17 ControlDecode.scala 72:17 ControlDecode.scala 79:17 ControlDecode.scala 85:17]
  assign io_memtoReg = io_rtype ? 1'h0 : _GEN_46; // @[ControlDecode.scala 29:17 ControlDecode.scala 49:17]
  assign io_memRead = io_rtype ? 1'h0 : _GEN_46; // @[ControlDecode.scala 30:17 ControlDecode.scala 50:17]
  assign io_memWrite = io_rtype ? 1'h0 : _GEN_47; // @[ControlDecode.scala 31:17 ControlDecode.scala 55:17]
  assign io_branch = io_rtype ? 1'h0 : _GEN_49; // @[ControlDecode.scala 32:17 ControlDecode.scala 61:17]
  assign io_oprndAsel = io_rtype ? 2'h0 : _GEN_51; // @[ControlDecode.scala 33:17 ControlDecode.scala 73:17 ControlDecode.scala 80:17 ControlDecode.scala 86:17]
  assign io_oprndBsel = io_rtype ? 1'h0 : _GEN_44; // @[ControlDecode.scala 34:17 ControlDecode.scala 44:17 ControlDecode.scala 51:17 ControlDecode.scala 56:17 ControlDecode.scala 67:17 ControlDecode.scala 74:17]
  assign io_immSel = io_rtype ? 2'h0 : _GEN_48; // @[ControlDecode.scala 35:17 ControlDecode.scala 57:17 ControlDecode.scala 68:17 ControlDecode.scala 75:17]
  assign io_nextPCsel = io_rtype ? 2'h0 : _GEN_50; // @[ControlDecode.scala 36:17 ControlDecode.scala 62:17 ControlDecode.scala 81:17 ControlDecode.scala 87:17]
  assign io_aluOP = io_rtype ? 3'h0 : _GEN_45; // @[ControlDecode.scala 37:17 ControlDecode.scala 45:17 ControlDecode.scala 52:17 ControlDecode.scala 58:17 ControlDecode.scala 63:17 ControlDecode.scala 69:17 ControlDecode.scala 76:17 ControlDecode.scala 82:17 ControlDecode.scala 88:17]
endmodule