module TypeDecode(
  input  [4:0] io_opcode,
  output       io_rtype,
  output       io_itype,
  output       io_load,
  output       io_stype,
  output       io_sbtype,
  output       io_lui,
  output       io_auipc,
  output       io_ujtype,
  output       io_jalr
);
  wire  _T; // @[TypeDecode.scala 29:22]
  wire  _T_1; // @[TypeDecode.scala 31:28]
  wire  _T_2; // @[TypeDecode.scala 33:28]
  wire  _T_3; // @[TypeDecode.scala 35:28]
  wire  _T_4; // @[TypeDecode.scala 37:28]
  wire  _T_5; // @[TypeDecode.scala 39:28]
  wire  _T_6; // @[TypeDecode.scala 41:28]
  wire  _T_7; // @[TypeDecode.scala 43:28]
  wire  _T_8; // @[TypeDecode.scala 45:28]
  wire  _GEN_2; // @[TypeDecode.scala 43:37]
  wire  _GEN_4; // @[TypeDecode.scala 41:37]
  wire  _GEN_5; // @[TypeDecode.scala 41:37]
  wire  _GEN_7; // @[TypeDecode.scala 39:37]
  wire  _GEN_8; // @[TypeDecode.scala 39:37]
  wire  _GEN_9; // @[TypeDecode.scala 39:37]
  wire  _GEN_11; // @[TypeDecode.scala 37:37]
  wire  _GEN_12; // @[TypeDecode.scala 37:37]
  wire  _GEN_13; // @[TypeDecode.scala 37:37]
  wire  _GEN_14; // @[TypeDecode.scala 37:37]
  wire  _GEN_16; // @[TypeDecode.scala 35:37]
  wire  _GEN_17; // @[TypeDecode.scala 35:37]
  wire  _GEN_18; // @[TypeDecode.scala 35:37]
  wire  _GEN_19; // @[TypeDecode.scala 35:37]
  wire  _GEN_20; // @[TypeDecode.scala 35:37]
  wire  _GEN_22; // @[TypeDecode.scala 33:37]
  wire  _GEN_23; // @[TypeDecode.scala 33:37]
  wire  _GEN_24; // @[TypeDecode.scala 33:37]
  wire  _GEN_25; // @[TypeDecode.scala 33:37]
  wire  _GEN_26; // @[TypeDecode.scala 33:37]
  wire  _GEN_27; // @[TypeDecode.scala 33:37]
  wire  _GEN_29; // @[TypeDecode.scala 31:37]
  wire  _GEN_30; // @[TypeDecode.scala 31:37]
  wire  _GEN_31; // @[TypeDecode.scala 31:37]
  wire  _GEN_32; // @[TypeDecode.scala 31:37]
  wire  _GEN_33; // @[TypeDecode.scala 31:37]
  wire  _GEN_34; // @[TypeDecode.scala 31:37]
  wire  _GEN_35; // @[TypeDecode.scala 31:37]
  assign _T = io_opcode == 5'hc; // @[TypeDecode.scala 29:22]
  assign _T_1 = io_opcode == 5'h4; // @[TypeDecode.scala 31:28]
  assign _T_2 = io_opcode == 5'h0; // @[TypeDecode.scala 33:28]
  assign _T_3 = io_opcode == 5'h8; // @[TypeDecode.scala 35:28]
  assign _T_4 = io_opcode == 5'h18; // @[TypeDecode.scala 37:28]
  assign _T_5 = io_opcode == 5'hd; // @[TypeDecode.scala 39:28]
  assign _T_6 = io_opcode == 5'h5; // @[TypeDecode.scala 41:28]
  assign _T_7 = io_opcode == 5'h1b; // @[TypeDecode.scala 43:28]
  assign _T_8 = io_opcode == 5'h19; // @[TypeDecode.scala 45:28]
  assign _GEN_2 = _T_7 ? 1'h0 : _T_8; // @[TypeDecode.scala 43:37]
  assign _GEN_4 = _T_6 ? 1'h0 : _T_7; // @[TypeDecode.scala 41:37]
  assign _GEN_5 = _T_6 ? 1'h0 : _GEN_2; // @[TypeDecode.scala 41:37]
  assign _GEN_7 = _T_5 ? 1'h0 : _T_6; // @[TypeDecode.scala 39:37]
  assign _GEN_8 = _T_5 ? 1'h0 : _GEN_4; // @[TypeDecode.scala 39:37]
  assign _GEN_9 = _T_5 ? 1'h0 : _GEN_5; // @[TypeDecode.scala 39:37]
  assign _GEN_11 = _T_4 ? 1'h0 : _T_5; // @[TypeDecode.scala 37:37]
  assign _GEN_12 = _T_4 ? 1'h0 : _GEN_7; // @[TypeDecode.scala 37:37]
  assign _GEN_13 = _T_4 ? 1'h0 : _GEN_8; // @[TypeDecode.scala 37:37]
  assign _GEN_14 = _T_4 ? 1'h0 : _GEN_9; // @[TypeDecode.scala 37:37]
  assign _GEN_16 = _T_3 ? 1'h0 : _T_4; // @[TypeDecode.scala 35:37]
  assign _GEN_17 = _T_3 ? 1'h0 : _GEN_11; // @[TypeDecode.scala 35:37]
  assign _GEN_18 = _T_3 ? 1'h0 : _GEN_12; // @[TypeDecode.scala 35:37]
  assign _GEN_19 = _T_3 ? 1'h0 : _GEN_13; // @[TypeDecode.scala 35:37]
  assign _GEN_20 = _T_3 ? 1'h0 : _GEN_14; // @[TypeDecode.scala 35:37]
  assign _GEN_22 = _T_2 ? 1'h0 : _T_3; // @[TypeDecode.scala 33:37]
  assign _GEN_23 = _T_2 ? 1'h0 : _GEN_16; // @[TypeDecode.scala 33:37]
  assign _GEN_24 = _T_2 ? 1'h0 : _GEN_17; // @[TypeDecode.scala 33:37]
  assign _GEN_25 = _T_2 ? 1'h0 : _GEN_18; // @[TypeDecode.scala 33:37]
  assign _GEN_26 = _T_2 ? 1'h0 : _GEN_19; // @[TypeDecode.scala 33:37]
  assign _GEN_27 = _T_2 ? 1'h0 : _GEN_20; // @[TypeDecode.scala 33:37]
  assign _GEN_29 = _T_1 ? 1'h0 : _T_2; // @[TypeDecode.scala 31:37]
  assign _GEN_30 = _T_1 ? 1'h0 : _GEN_22; // @[TypeDecode.scala 31:37]
  assign _GEN_31 = _T_1 ? 1'h0 : _GEN_23; // @[TypeDecode.scala 31:37]
  assign _GEN_32 = _T_1 ? 1'h0 : _GEN_24; // @[TypeDecode.scala 31:37]
  assign _GEN_33 = _T_1 ? 1'h0 : _GEN_25; // @[TypeDecode.scala 31:37]
  assign _GEN_34 = _T_1 ? 1'h0 : _GEN_26; // @[TypeDecode.scala 31:37]
  assign _GEN_35 = _T_1 ? 1'h0 : _GEN_27; // @[TypeDecode.scala 31:37]
  assign io_rtype = io_opcode == 5'hc; // @[TypeDecode.scala 19:19 TypeDecode.scala 30:19]
  assign io_itype = _T ? 1'h0 : _T_1; // @[TypeDecode.scala 20:19 TypeDecode.scala 32:19]
  assign io_load = _T ? 1'h0 : _GEN_29; // @[TypeDecode.scala 21:19 TypeDecode.scala 34:19]
  assign io_stype = _T ? 1'h0 : _GEN_30; // @[TypeDecode.scala 22:19 TypeDecode.scala 36:19]
  assign io_sbtype = _T ? 1'h0 : _GEN_31; // @[TypeDecode.scala 23:19 TypeDecode.scala 38:19]
  assign io_lui = _T ? 1'h0 : _GEN_32; // @[TypeDecode.scala 24:19 TypeDecode.scala 40:19]
  assign io_auipc = _T ? 1'h0 : _GEN_33; // @[TypeDecode.scala 25:19 TypeDecode.scala 42:19]
  assign io_ujtype = _T ? 1'h0 : _GEN_34; // @[TypeDecode.scala 26:19 TypeDecode.scala 44:19]
  assign io_jalr = _T ? 1'h0 : _GEN_35; // @[TypeDecode.scala 27:19 TypeDecode.scala 46:19]
endmodule